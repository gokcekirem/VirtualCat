library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity HUDREDHZ_CLOCK_GENERATOR is
    Port ( MCLK : in  STD_LOGIC;
           HUNDREDHZCLOCK : out  STD_LOGIC);
end HUDREDHZ_CLOCK_GENERATOR;

architecture Behavioral of HUDREDHZ_CLOCK_GENERATOR is

SIGNAL COUNTER : STD_LOGIC_VECTOR(20 DOWNTO 0) := "000000000000000000000";

begin

CLK_PROCESS: PROCESS(MCLK)

BEGIN
	--INCREMENT COUNTER
	IF(MCLK'EVENT AND MCLK = '1') THEN
		IF(COUNTER < "111101000010010000000") THEN 
			COUNTER <= COUNTER + "110"; 
		ELSE
			COUNTER <= "000000000000000000000";
		END IF;	
	END IF;
END PROCESS;
--END OF CLOCK PROCESS

HUNDREDHZCLOCK <= '1' WHEN COUNTER < "011110100001001000000" ELSE '0';

end Behavioral;

