
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

ENTITY SSSLIB IS
    PORT ( 
				MCLK							: IN  STD_LOGIC;
				B1,B2,B3,B4		 		   : IN STD_LOGIC;
				SW0,SW1,SW2					: IN STD_LOGIC;
				SEVSEG_DATA					: OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
            SEVSEG_CONTROL				: OUT  STD_LOGIC_VECTOR (7 DOWNTO 0));
END SSSLIB;

ARCHITECTURE BEHAVIORAL OF SSSLIB IS

--INTERMEDIATE SIGNALS
SIGNAL WIRE_HUNDREDHZ_CLOCK : STD_LOGIC;
SIGNAL WIRE_oneHZ_CLOCK : STD_LOGIC;

SIGNAL WIRE_SEVSEG_DATA		 : STD_LOGIC_VECTOR(4 DOWNTO 0);

SIGNAL WIRE_SEVSEG_DRIVER :STD_LOGIC_VECTOR(7 DOWNTO 0);


BEGIN

--ADD CLOCK GENERATOR
CLOCK_GENERATOR : ENTITY WORK.HUDREDHZ_CLOCK_GENERATOR PORT MAP(
	MCLK => MCLK,
	HUNDREDHZCLOCK => WIRE_HUNDREDHZ_CLOCK
		
	
);

--ADD DRIVER
CAT : ENTITY WORK.CAT PORT MAP(
 oneHZCLOCK => WIRE_oneHZ_CLOCK,
 
 B1 => B1,
 B2 => B2,
 B3 => B3,
 B4 => B4,
 sw0 		=> sw0,
 sw1 		=> sw1,
 sw2 		=> sw2,

 CLK => WIRE_HUNDREDHZ_CLOCK,
 
 SEV_SEG_DATA => WIRE_SEVSEG_DATA,
 SEV_SEG_DRIVER => WIRE_SEVSEG_DRIVER
);

oneHZ_CLOCK: ENTITY WORK.oneHZ_CLOCK_GENERATOR PORT MAP(
 mclk => mclk,
 oneHZCLOCK  => WIRE_oneHZ_CLOCK
 
);

--ADD DECODER
DECODER : ENTITY WORK.SEVSEG_DECODER PORT MAP(

	SEV_SEG_DATA => WIRE_SEVSEG_DATA,
	 SEV_SEG_DRIVER => WIRE_SEVSEG_DRIVER,

	SEVSEG_BUS => SEVSEG_DATA,
	
	 SEVSEG_CONTROL  => SEVSEG_CONTROL 
	
	
	);

END BEHAVIORAL;

